interface spi_if;
  logic clk;
  logic rst;
  logic newdata;
  logic [11:0] din;
  logic sclk;
  logic cs;
  logic mosi;
  
endinterface
